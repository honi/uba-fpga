library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package stopwatch_pkg is
    type matrix is array (integer range <>) of std_logic_vector(3 downto 0);
end package;
